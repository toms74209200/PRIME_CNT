-- =====================================================================
--  Title       : Prime number counter
--
--  File Name	: PRIME_CNT.vhd
--  Project     :
--  Block       :
--  Tree        :
--  Designer    : toms74209200 <https://github.com/toms74209200>
--  Created     : 2019/03/14
--  Copyright   : 2019 toms74209200
--  License     : MIT License.
--                http://opensource.org/licenses/mit-license.php
-- =====================================================================
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity PRIME_CNT is
    port(
    -- System --
        CLK     : in    std_logic;                      --(p) Clock
        nRST    : in    std_logic;                      --(n) Reset

    -- Control --
        STR     : in    std_logic;                      --(p) Start pulse
        BUSY    : out   std_logic;                      --(p) Calculation busy
        VALID   : out   std_logic;                      --(p) Data valid

    -- Data --
        DAT     : out	std_logic_vector(31 downto 0)   --(p) Data
        );
end PRIME_CNT;

architecture RTL of PRIME_CNT is

-- Parameter --
constant CalcMax        : std_logic_vector(31 downto 0) := X"05F5_E0FF";    -- Calculation max 99,999,999
constant PrimeMax       : integer := 1227;                                  -- ROM max prime order

-- Internal signals --
signal busy_i           : std_logic;                        --(p) Calculation busy
signal valid_i          : std_logic;                        --(p) Data valid
signal dat_i            : std_logic_vector(DAT'range);      --(p) Data
signal cnt_pls          : std_logic_vector(0 to PrimeMax);  --(p) Prime counter pulse

-- Data array --
type PrimeDatType       is array(0 to 1227) of std_logic_vector(15 downto 0);
signal ary_prime_cnt    : PrimeDatType;

-- ROM table --
constant rom_prime      : PrimeDatType :=
(
    X"0003",
    X"0005",
    X"0007",
    X"000B",
    X"000D",
    X"0011",
    X"0013",
    X"0017",
    X"001D",
    X"001F",
    X"0025",
    X"0029",
    X"002B",
    X"002F",
    X"0035",
    X"003B",
    X"003D",
    X"0043",
    X"0047",
    X"0049",
    X"004F",
    X"0053",
    X"0059",
    X"0061",
    X"0065",
    X"0067",
    X"006B",
    X"006D",
    X"0071",
    X"007F",
    X"0083",
    X"0089",
    X"008B",
    X"0095",
    X"0097",
    X"009D",
    X"00A3",
    X"00A7",
    X"00AD",
    X"00B3",
    X"00B5",
    X"00BF",
    X"00C1",
    X"00C5",
    X"00C7",
    X"00D3",
    X"00DF",
    X"00E3",
    X"00E5",
    X"00E9",
    X"00EF",
    X"00F1",
    X"00FB",
    X"0101",
    X"0107",
    X"010D",
    X"010F",
    X"0115",
    X"0119",
    X"011B",
    X"0125",
    X"0133",
    X"0137",
    X"0139",
    X"013D",
    X"014B",
    X"0151",
    X"015B",
    X"015D",
    X"0161",
    X"0167",
    X"016F",
    X"0175",
    X"017B",
    X"017F",
    X"0185",
    X"018D",
    X"0191",
    X"0199",
    X"01A3",
    X"01A5",
    X"01AF",
    X"01B1",
    X"01B7",
    X"01BB",
    X"01C1",
    X"01C9",
    X"01CD",
    X"01CF",
    X"01D3",
    X"01DF",
    X"01E7",
    X"01EB",
    X"01F3",
    X"01F7",
    X"01FD",
    X"0209",
    X"020B",
    X"021D",
    X"0223",
    X"022D",
    X"0233",
    X"0239",
    X"023B",
    X"0241",
    X"024B",
    X"0251",
    X"0257",
    X"0259",
    X"025F",
    X"0265",
    X"0269",
    X"026B",
    X"0277",
    X"0281",
    X"0283",
    X"0287",
    X"028D",
    X"0293",
    X"0295",
    X"02A1",
    X"02A5",
    X"02AB",
    X"02B3",
    X"02BD",
    X"02C5",
    X"02CF",
    X"02D7",
    X"02DD",
    X"02E3",
    X"02E7",
    X"02EF",
    X"02F5",
    X"02F9",
    X"0301",
    X"0305",
    X"0313",
    X"031D",
    X"0329",
    X"032B",
    X"0335",
    X"0337",
    X"033B",
    X"033D",
    X"0347",
    X"0355",
    X"0359",
    X"035B",
    X"035F",
    X"036D",
    X"0371",
    X"0373",
    X"0377",
    X"038B",
    X"038F",
    X"0397",
    X"03A1",
    X"03A9",
    X"03AD",
    X"03B3",
    X"03B9",
    X"03C7",
    X"03CB",
    X"03D1",
    X"03D7",
    X"03DF",
    X"03E5",
    X"03F1",
    X"03F5",
    X"03FB",
    X"03FD",
    X"0407",
    X"0409",
    X"040F",
    X"0419",
    X"041B",
    X"0425",
    X"0427",
    X"042D",
    X"043F",
    X"0443",
    X"0445",
    X"0449",
    X"044F",
    X"0455",
    X"045D",
    X"0463",
    X"0469",
    X"047F",
    X"0481",
    X"048B",
    X"0493",
    X"049D",
    X"04A3",
    X"04A9",
    X"04B1",
    X"04BD",
    X"04C1",
    X"04C7",
    X"04CD",
    X"04CF",
    X"04D5",
    X"04E1",
    X"04EB",
    X"04FD",
    X"04FF",
    X"0503",
    X"0509",
    X"050B",
    X"0511",
    X"0515",
    X"0517",
    X"051B",
    X"0527",
    X"0529",
    X"052F",
    X"0551",
    X"0557",
    X"055D",
    X"0565",
    X"0577",
    X"0581",
    X"058F",
    X"0593",
    X"0595",
    X"0599",
    X"059F",
    X"05A7",
    X"05AB",
    X"05AD",
    X"05B3",
    X"05BF",
    X"05C9",
    X"05CB",
    X"05CF",
    X"05D1",
    X"05D5",
    X"05DB",
    X"05E7",
    X"05F3",
    X"05FB",
    X"0607",
    X"060D",
    X"0611",
    X"0617",
    X"061F",
    X"0623",
    X"062B",
    X"062F",
    X"063D",
    X"0641",
    X"0647",
    X"0649",
    X"064D",
    X"0653",
    X"0655",
    X"065B",
    X"0665",
    X"0679",
    X"067F",
    X"0683",
    X"0685",
    X"069D",
    X"06A1",
    X"06A3",
    X"06AD",
    X"06B9",
    X"06BB",
    X"06C5",
    X"06CD",
    X"06D3",
    X"06D9",
    X"06DF",
    X"06F1",
    X"06F7",
    X"06FB",
    X"06FD",
    X"0709",
    X"0713",
    X"071F",
    X"0727",
    X"0737",
    X"0745",
    X"074B",
    X"074F",
    X"0751",
    X"0755",
    X"0757",
    X"0761",
    X"076D",
    X"0773",
    X"0779",
    X"078B",
    X"078D",
    X"079D",
    X"079F",
    X"07B5",
    X"07BB",
    X"07C3",
    X"07C9",
    X"07CD",
    X"07CF",
    X"07D3",
    X"07DB",
    X"07E1",
    X"07EB",
    X"07ED",
    X"07F7",
    X"0805",
    X"080F",
    X"0815",
    X"0821",
    X"0823",
    X"0827",
    X"0829",
    X"0833",
    X"083F",
    X"0841",
    X"0851",
    X"0853",
    X"0859",
    X"085D",
    X"085F",
    X"0869",
    X"0871",
    X"0883",
    X"089B",
    X"089F",
    X"08A5",
    X"08AD",
    X"08BD",
    X"08BF",
    X"08C3",
    X"08CB",
    X"08DB",
    X"08DD",
    X"08E1",
    X"08E9",
    X"08EF",
    X"08F5",
    X"08F9",
    X"0905",
    X"0907",
    X"091D",
    X"0923",
    X"0925",
    X"092B",
    X"092F",
    X"0935",
    X"0943",
    X"0949",
    X"094D",
    X"094F",
    X"0955",
    X"0959",
    X"095F",
    X"096B",
    X"0971",
    X"0977",
    X"0985",
    X"0989",
    X"098F",
    X"099B",
    X"09A3",
    X"09A9",
    X"09AD",
    X"09C7",
    X"09D9",
    X"09E3",
    X"09EB",
    X"09EF",
    X"09F5",
    X"09F7",
    X"09FD",
    X"0A13",
    X"0A1F",
    X"0A21",
    X"0A31",
    X"0A39",
    X"0A3D",
    X"0A49",
    X"0A57",
    X"0A61",
    X"0A63",
    X"0A67",
    X"0A6F",
    X"0A75",
    X"0A7B",
    X"0A7F",
    X"0A81",
    X"0A85",
    X"0A8B",
    X"0A93",
    X"0A97",
    X"0A99",
    X"0A9F",
    X"0AA9",
    X"0AAB",
    X"0AB5",
    X"0ABD",
    X"0AC1",
    X"0ACF",
    X"0AD9",
    X"0AE5",
    X"0AE7",
    X"0AED",
    X"0AF1",
    X"0AF3",
    X"0B03",
    X"0B11",
    X"0B15",
    X"0B1B",
    X"0B23",
    X"0B29",
    X"0B2D",
    X"0B3F",
    X"0B47",
    X"0B51",
    X"0B57",
    X"0B5D",
    X"0B65",
    X"0B6F",
    X"0B7B",
    X"0B89",
    X"0B8D",
    X"0B93",
    X"0B99",
    X"0B9B",
    X"0BB7",
    X"0BB9",
    X"0BC3",
    X"0BCB",
    X"0BCF",
    X"0BDD",
    X"0BE1",
    X"0BE9",
    X"0BF5",
    X"0BFB",
    X"0C07",
    X"0C0B",
    X"0C11",
    X"0C25",
    X"0C2F",
    X"0C31",
    X"0C41",
    X"0C5B",
    X"0C5F",
    X"0C61",
    X"0C6D",
    X"0C73",
    X"0C77",
    X"0C83",
    X"0C89",
    X"0C91",
    X"0C95",
    X"0C9D",
    X"0CB3",
    X"0CB5",
    X"0CB9",
    X"0CBB",
    X"0CC7",
    X"0CE3",
    X"0CE5",
    X"0CEB",
    X"0CF1",
    X"0CF7",
    X"0CFB",
    X"0D01",
    X"0D03",
    X"0D0F",
    X"0D13",
    X"0D1F",
    X"0D21",
    X"0D2B",
    X"0D2D",
    X"0D3D",
    X"0D3F",
    X"0D4F",
    X"0D55",
    X"0D69",
    X"0D79",
    X"0D81",
    X"0D85",
    X"0D87",
    X"0D8B",
    X"0D8D",
    X"0DA3",
    X"0DAB",
    X"0DB7",
    X"0DBD",
    X"0DC7",
    X"0DC9",
    X"0DCD",
    X"0DD3",
    X"0DD5",
    X"0DDB",
    X"0DE5",
    X"0DE7",
    X"0DF3",
    X"0DFD",
    X"0DFF",
    X"0E09",
    X"0E17",
    X"0E1D",
    X"0E21",
    X"0E27",
    X"0E2F",
    X"0E35",
    X"0E3B",
    X"0E4B",
    X"0E57",
    X"0E59",
    X"0E5D",
    X"0E6B",
    X"0E71",
    X"0E75",
    X"0E7D",
    X"0E87",
    X"0E8F",
    X"0E95",
    X"0E9B",
    X"0EB1",
    X"0EB7",
    X"0EB9",
    X"0EC3",
    X"0ED1",
    X"0ED5",
    X"0EDB",
    X"0EED",
    X"0EEF",
    X"0EF9",
    X"0F07",
    X"0F0B",
    X"0F0D",
    X"0F17",
    X"0F25",
    X"0F29",
    X"0F31",
    X"0F43",
    X"0F47",
    X"0F4D",
    X"0F4F",
    X"0F53",
    X"0F59",
    X"0F5B",
    X"0F67",
    X"0F6B",
    X"0F7F",
    X"0F95",
    X"0FA1",
    X"0FA3",
    X"0FA7",
    X"0FAD",
    X"0FB3",
    X"0FB5",
    X"0FBB",
    X"0FD1",
    X"0FD3",
    X"0FD9",
    X"0FE9",
    X"0FEF",
    X"0FFB",
    X"0FFD",
    X"1003",
    X"100F",
    X"101F",
    X"1021",
    X"1025",
    X"102B",
    X"1039",
    X"103D",
    X"103F",
    X"1051",
    X"1069",
    X"1073",
    X"1079",
    X"107B",
    X"1085",
    X"1087",
    X"1091",
    X"1093",
    X"109D",
    X"10A3",
    X"10A5",
    X"10AF",
    X"10B1",
    X"10BB",
    X"10C1",
    X"10C9",
    X"10E7",
    X"10F1",
    X"10F3",
    X"10FD",
    X"1105",
    X"110B",
    X"1115",
    X"1127",
    X"112D",
    X"1139",
    X"1145",
    X"1147",
    X"1159",
    X"115F",
    X"1163",
    X"1169",
    X"116F",
    X"1181",
    X"1183",
    X"118D",
    X"119B",
    X"11A1",
    X"11A5",
    X"11A7",
    X"11AB",
    X"11C3",
    X"11C5",
    X"11D1",
    X"11D7",
    X"11E7",
    X"11EF",
    X"11F5",
    X"11FB",
    X"120D",
    X"121D",
    X"121F",
    X"1223",
    X"1229",
    X"122B",
    X"1231",
    X"1237",
    X"1241",
    X"1247",
    X"1253",
    X"125F",
    X"1271",
    X"1273",
    X"1279",
    X"127D",
    X"128F",
    X"1297",
    X"12AF",
    X"12B3",
    X"12B5",
    X"12B9",
    X"12BF",
    X"12C1",
    X"12CD",
    X"12D1",
    X"12DF",
    X"12FD",
    X"1307",
    X"130D",
    X"1319",
    X"1327",
    X"132D",
    X"1337",
    X"1343",
    X"1345",
    X"1349",
    X"134F",
    X"1357",
    X"135D",
    X"1367",
    X"1369",
    X"136D",
    X"137B",
    X"1381",
    X"1387",
    X"138B",
    X"1391",
    X"1393",
    X"139D",
    X"139F",
    X"13AF",
    X"13BB",
    X"13C3",
    X"13D5",
    X"13D9",
    X"13DF",
    X"13EB",
    X"13ED",
    X"13F3",
    X"13F9",
    X"13FF",
    X"141B",
    X"1421",
    X"142F",
    X"1433",
    X"143B",
    X"1445",
    X"144D",
    X"1459",
    X"146B",
    X"146F",
    X"1471",
    X"1475",
    X"148D",
    X"1499",
    X"149F",
    X"14A1",
    X"14B1",
    X"14B7",
    X"14BD",
    X"14CB",
    X"14D5",
    X"14E3",
    X"14E7",
    X"1505",
    X"150B",
    X"1511",
    X"1517",
    X"151F",
    X"1525",
    X"1529",
    X"152B",
    X"1537",
    X"153D",
    X"1541",
    X"1543",
    X"1549",
    X"155F",
    X"1565",
    X"1567",
    X"156B",
    X"157D",
    X"157F",
    X"1583",
    X"158F",
    X"1591",
    X"1597",
    X"159B",
    X"15B5",
    X"15BB",
    X"15C1",
    X"15C5",
    X"15CD",
    X"15D7",
    X"15F7",
    X"1607",
    X"1609",
    X"160F",
    X"1613",
    X"1615",
    X"1619",
    X"161B",
    X"1625",
    X"1633",
    X"1639",
    X"163D",
    X"1645",
    X"164F",
    X"1655",
    X"1669",
    X"166D",
    X"166F",
    X"1675",
    X"1693",
    X"1697",
    X"169F",
    X"16A9",
    X"16AF",
    X"16B5",
    X"16BD",
    X"16C3",
    X"16CF",
    X"16D3",
    X"16D9",
    X"16DB",
    X"16E1",
    X"16E5",
    X"16EB",
    X"16ED",
    X"16F7",
    X"16F9",
    X"1709",
    X"170F",
    X"1723",
    X"1727",
    X"1733",
    X"1741",
    X"175D",
    X"1763",
    X"1777",
    X"177B",
    X"178D",
    X"1795",
    X"179B",
    X"179F",
    X"17A5",
    X"17B3",
    X"17B9",
    X"17BF",
    X"17C9",
    X"17CB",
    X"17D5",
    X"17E1",
    X"17E9",
    X"17F3",
    X"17F5",
    X"17FF",
    X"1807",
    X"1813",
    X"181D",
    X"1835",
    X"1837",
    X"183B",
    X"1843",
    X"1849",
    X"184D",
    X"1855",
    X"1867",
    X"1871",
    X"1877",
    X"187D",
    X"187F",
    X"1885",
    X"188F",
    X"189B",
    X"189D",
    X"18A7",
    X"18AD",
    X"18B3",
    X"18B9",
    X"18C1",
    X"18C7",
    X"18D1",
    X"18D7",
    X"18D9",
    X"18DF",
    X"18E5",
    X"18EB",
    X"18F5",
    X"18FD",
    X"1915",
    X"191B",
    X"1931",
    X"1933",
    X"1945",
    X"1949",
    X"1951",
    X"195B",
    X"1979",
    X"1981",
    X"1993",
    X"1997",
    X"1999",
    X"19A3",
    X"19A9",
    X"19AB",
    X"19B1",
    X"19B5",
    X"19C7",
    X"19CF",
    X"19DB",
    X"19ED",
    X"19FD",
    X"1A03",
    X"1A05",
    X"1A11",
    X"1A17",
    X"1A21",
    X"1A23",
    X"1A2D",
    X"1A2F",
    X"1A35",
    X"1A3F",
    X"1A4D",
    X"1A51",
    X"1A69",
    X"1A6B",
    X"1A7B",
    X"1A7D",
    X"1A87",
    X"1A89",
    X"1A93",
    X"1AA7",
    X"1AAB",
    X"1AAD",
    X"1AB1",
    X"1AB9",
    X"1AC9",
    X"1ACF",
    X"1AD5",
    X"1AD7",
    X"1AE3",
    X"1AF3",
    X"1AFB",
    X"1AFF",
    X"1B05",
    X"1B23",
    X"1B25",
    X"1B2F",
    X"1B31",
    X"1B37",
    X"1B3B",
    X"1B41",
    X"1B47",
    X"1B4F",
    X"1B55",
    X"1B59",
    X"1B65",
    X"1B6B",
    X"1B73",
    X"1B7F",
    X"1B83",
    X"1B91",
    X"1B9D",
    X"1BA7",
    X"1BBF",
    X"1BC5",
    X"1BD1",
    X"1BD7",
    X"1BD9",
    X"1BEF",
    X"1BF7",
    X"1C09",
    X"1C13",
    X"1C19",
    X"1C27",
    X"1C2B",
    X"1C2D",
    X"1C33",
    X"1C3D",
    X"1C45",
    X"1C4B",
    X"1C4F",
    X"1C55",
    X"1C73",
    X"1C81",
    X"1C8B",
    X"1C8D",
    X"1C99",
    X"1CA3",
    X"1CA5",
    X"1CB5",
    X"1CB7",
    X"1CC9",
    X"1CE1",
    X"1CF3",
    X"1CF9",
    X"1D09",
    X"1D1B",
    X"1D21",
    X"1D23",
    X"1D35",
    X"1D39",
    X"1D3F",
    X"1D41",
    X"1D4B",
    X"1D53",
    X"1D5D",
    X"1D63",
    X"1D69",
    X"1D71",
    X"1D75",
    X"1D7B",
    X"1D7D",
    X"1D87",
    X"1D89",
    X"1D95",
    X"1D99",
    X"1D9F",
    X"1DA5",
    X"1DA7",
    X"1DB3",
    X"1DB7",
    X"1DC5",
    X"1DD7",
    X"1DDB",
    X"1DE1",
    X"1DF5",
    X"1DF9",
    X"1E01",
    X"1E07",
    X"1E0B",
    X"1E13",
    X"1E17",
    X"1E25",
    X"1E2B",
    X"1E2F",
    X"1E3D",
    X"1E49",
    X"1E4D",
    X"1E4F",
    X"1E6D",
    X"1E71",
    X"1E89",
    X"1E8F",
    X"1E95",
    X"1EA1",
    X"1EAD",
    X"1EBB",
    X"1EC1",
    X"1EC5",
    X"1EC7",
    X"1ECB",
    X"1EDD",
    X"1EE3",
    X"1EEF",
    X"1EF7",
    X"1EFD",
    X"1F01",
    X"1F0D",
    X"1F0F",
    X"1F1B",
    X"1F39",
    X"1F49",
    X"1F4B",
    X"1F51",
    X"1F67",
    X"1F75",
    X"1F7B",
    X"1F85",
    X"1F91",
    X"1F97",
    X"1F99",
    X"1F9D",
    X"1FA5",
    X"1FAF",
    X"1FB5",
    X"1FBB",
    X"1FD3",
    X"1FE1",
    X"1FE7",
    X"1FEB",
    X"1FF3",
    X"1FFF",
    X"2011",
    X"201B",
    X"201D",
    X"2027",
    X"2029",
    X"202D",
    X"2033",
    X"2047",
    X"204D",
    X"2051",
    X"205F",
    X"2063",
    X"2065",
    X"2069",
    X"2077",
    X"207D",
    X"2089",
    X"20A1",
    X"20AB",
    X"20B1",
    X"20B9",
    X"20C3",
    X"20C5",
    X"20E3",
    X"20E7",
    X"20ED",
    X"20EF",
    X"20FB",
    X"20FF",
    X"210D",
    X"2113",
    X"2135",
    X"2141",
    X"2149",
    X"214F",
    X"2159",
    X"215B",
    X"215F",
    X"2173",
    X"217D",
    X"2185",
    X"2195",
    X"2197",
    X"21A1",
    X"21AF",
    X"21B3",
    X"21B5",
    X"21C1",
    X"21C7",
    X"21D7",
    X"21DD",
    X"21E5",
    X"21E9",
    X"21F1",
    X"21F5",
    X"21FB",
    X"2203",
    X"2209",
    X"220F",
    X"221B",
    X"2221",
    X"2225",
    X"222B",
    X"2231",
    X"2239",
    X"224B",
    X"224F",
    X"2263",
    X"2267",
    X"2273",
    X"2275",
    X"227F",
    X"2285",
    X"2287",
    X"2291",
    X"229D",
    X"229F",
    X"22A3",
    X"22B7",
    X"22BD",
    X"22DB",
    X"22E1",
    X"22E5",
    X"22ED",
    X"22F7",
    X"2303",
    X"2309",
    X"230B",
    X"2327",
    X"2329",
    X"232F",
    X"2333",
    X"2335",
    X"2345",
    X"2351",
    X"2353",
    X"2359",
    X"2363",
    X"236B",
    X"2383",
    X"238F",
    X"2395",
    X"23A7",
    X"23AD",
    X"23B1",
    X"23BF",
    X"23C5",
    X"23C9",
    X"23D5",
    X"23DD",
    X"23E3",
    X"23EF",
    X"23F3",
    X"23F9",
    X"2405",
    X"240B",
    X"2417",
    X"2419",
    X"2429",
    X"243D",
    X"2441",
    X"2443",
    X"244D",
    X"245F",
    X"2467",
    X"246B",
    X"2479",
    X"247D",
    X"247F",
    X"2485",
    X"249B",
    X"24A1",
    X"24AF",
    X"24B5",
    X"24BB",
    X"24C5",
    X"24CB",
    X"24CD",
    X"24D7",
    X"24D9",
    X"24DD",
    X"24DF",
    X"24F5",
    X"24F7",
    X"24FB",
    X"2501",
    X"2507",
    X"2513",
    X"2519",
    X"2527",
    X"2531",
    X"253D",
    X"2543",
    X"254B",
    X"254F",
    X"2573",
    X"2581",
    X"258D",
    X"2593",
    X"2597",
    X"259D",
    X"259F",
    X"25AB",
    X"25B1",
    X"25BD",
    X"25CD",
    X"25CF",
    X"25D9",
    X"25E1",
    X"25F7",
    X"25F9",
    X"2605",
    X"260B",
    X"260F",
    X"2615",
    X"2627",
    X"2629",
    X"2635",
    X"263B",
    X"263F",
    X"264B",
    X"2653",
    X"2659",
    X"2665",
    X"2669",
    X"266F",
    X"267B",
    X"2681",
    X"2683",
    X"268F",
    X"269B",
    X"269F",
    X"26AD",
    X"26B3",
    X"26C3",
    X"26C9",
    X"26CB",
    X"26D5",
    X"26DD",
    X"26EF",
    X"26F5"
);

begin
-- ***********************************************************
--  Busy flag
-- ***********************************************************
process (CLK, nRST) begin
    if (nRST = '0') then
        busy_i <= '0';
    elsif (CLK'event and CLK = '1') then
        if (dat_i = CalcMax) then
            busy_i <= '0';
        elsif (STR = '1') then
            busy_i <= '1';
        end if;
    end if;
end process;

BUSY <= busy_i;


-- ***********************************************************
--  Prime number counter
-- ***********************************************************
process (CLK, nRST) begin
    for i in cnt_pls'range loop
        if (nRST = '0') then
            ary_prime_cnt(i) <= (others => '0');
        elsif (CLK'event and CLK = '1') then
            if (busy_i = '1') then
                if (dat_i = rom_prime(i)) then
                    ary_prime_cnt(i) <= rom_prime(i);
                elsif (ary_prime_cnt(i) = rom_prime(i)) then
                    ary_prime_cnt(i) <= X"0001";
                else
                    ary_prime_cnt(i) <= ary_prime_cnt(i) + 1;
                end if;
            else
                ary_prime_cnt(i) <= (others => '0');
            end if;
        end if;
    end loop;
end process;

ARY_CNT_PLS : for i in cnt_pls'range generate
    cnt_pls(i) <= '1' when (ary_prime_cnt(i) = rom_prime(i)-1) else '0';
end generate;


-- ***********************************************************
--  Data counter
-- ***********************************************************
process (CLK, nRST) begin
    if (nRST = '0') then
        dat_i <= (others => '0');
    elsif (CLK'event and CLK = '1') then
        if (busy_i = '1') then
            if (dat_i = CalcMax) then
                dat_i <= X"0000_0001";
            else
                dat_i <= dat_i + 2;
            end if;
        else
            dat_i <= X"0000_0001";
        end if;
    end if;
end process;


-- ***********************************************************
--  Data
-- ***********************************************************
DAT <= dat_i when (valid_i = '1') else (others => '0');


-- ***********************************************************
--  Data valid
-- ***********************************************************
valid_i <= '1' when (busy_i = '1' and cnt_pls = 0) else '0';

VALID <= valid_i;


end RTL; --PRIME_CNT